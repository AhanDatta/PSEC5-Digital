// Interface with DUT to the rest of the system, includes all inputs and outputs
interface intf(input logic clk);

  logic rstn;
  logic iclk;
  logic sclk;
  logic ch0;
  logic ch1;
  logic ch2;
  logic ch3;
  logic ch4;
  logic ch5;
  logic ch6;
  logic ch7;
  logic serial_in;
  logic serial_out;

//***NEED TO INCLUDE CLOCKING BLOCKS AND MODPORTS!!!


endinterface